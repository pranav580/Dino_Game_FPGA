module Huddle(
	clk,
	rst,
	breakGameFlag,
	hor_reg,
	ver_reg,
	hudPosHorFrom,hudPosHorTo,hudPosVerFrom,hudPosVerTo
);

input clk,rst,hor_reg,ver_reg,breakGameFlag;
output reg hudPosHorFrom,hudPosHorTo,hudPosVerFrom,hudPosVerTo;


endmodule
