module Score(clk,rst,BreakFlag,scoreHorFrom,scoreHorTo,scoreVerFrom,scoreVerTo);

input clk,rst,BreakFlag;
output reg scoreHorFrom,scoreHorTo,scoreVerFrom,scoreVerTo;



endmodule
