module Score(clk,rst,BreakFlag,scoreHorFrom,scoreHorTo,scoreVerFrom,scoreVerTo);

input clk,rst,BreakFlag;
output reg scoreHorFrom,scoreHorTo,scoreVerFrom,scoreVerTE:\Bhavesh\SVVV_DOCS\FPGA\Dino_Game_(3)\Dino_Game_FPGA>;



endmodule
